library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity stage1_twiddle_i_rom is
    generic (
        ADDR_WIDTH : POSITIVE := 6;
        DATA_WIDTH : POSITIVE := 16
    );
    port (
        addr : in std_logic_vector(ADDR_WIDTH - 1 downto 0);
        dout : out std_logic_vector(DATA_WIDTH - 1 downto 0)
    );
end;
architecture rtl of stage1_twiddle_i_rom is
    type mem_type is array (0 to (2 ** ADDR_WIDTH) - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);
    constant memory : mem_type := ("0000000000000000", "1111001110000100", "1110011110000010", "1101110001110010", "1101001010111111", "1100101011001001", "1100010011011111", "1100000100111011", "1100000000000000", "1100000100111011", "1100010011011111", "1100101011001001", "1101001010111111", "1101110001110010", "1110011110000010", "1111001110000100", "0000000000000000", "1111100110111010", "1111001110000100", "1110110101101100", "1110011110000010", "1110000111010101", "1101110001110010", "1101011101100110", "1101001010111111", "1100111010000111", "1100101011001001", "1100011110001111", "1100010011011111", "1100001011000001", "1100000100111011", "1100000001001111", "0000000000000000", "1110110101101100", "1101110001110010", "1100111010000111", "1100010011011111", "1100000001001111", "1100000100111011", "1100011110001111", "1101001010111111", "1110000111010101", "1111001110000100", "0000011001000110", "0001100001111110", "0010100010011010", "0011010100110111", "0011110100111111", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000", "0000000000000000");
begin
    dout <= std_logic_vector(memory(CONV_INTEGER(addr)));
end;
